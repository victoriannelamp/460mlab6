module bcd(); 

endmodule 