module tracker(); 

endmodule 