module pulse_gen_clk_div(clk,rst,start,mode, pusle, clk_60hz); 
input clk,rst, start, mode; 
output pulse,clk_60hz; 

endmodule 